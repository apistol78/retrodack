input CLOCK,
output LCD_VSYNC,
output LCD_HSYNC,
output LCD_B0,
output LCD_G2,
output LCD_G3,
output LCD_G5,
output LCD_CS,
output LCD_R3,
output LCD_R2,
output LCD_R4,
output LCD_R5,
output LCD_B5,
output LCD_B4,
output LCD_B3,
output LCD_CLK,
output LCD_ENABLE,
output LCD_B1,
output LCD_B2,
output LCD_G0,
output LCD_G1,
output LCD_G4,
output LCD_BACKLIGHT_CTRL,
output LCD_R0,
output LCD_R1,
output UART_TX,
input UART_RX,
inout SD_DAT1,
inout SD_DAT0,
output SD_CLK,
output SD_CMD,
inout SD_DAT3,
inout SD_DAT2,
input USE_HCI_INT,
output USE_HCI_MOSI,
input USE_HCI_MISO,
output USE_HCI_SS_n,
output USE_HCI_SCLK,
output USB_HCI_RESET_n
