input CLOCK,
output LED_G,
output LED_R,
output LED_B,
output LCD_VSYNC,
output LCD_HSYNC,
output LCD_B0,
output LCD_G2,
output LCD_G3,
output LCD_G5,
output LCD_CS,
output LCD_R3,
output LCD_R2,
output LCD_R4,
output LCD_R5,
output LCD_B5,
output LCD_B4,
output LCD_B3,
output LCD_CLK,
output LCD_ENABLE,
output LCD_B1,
output LCD_B2,
output LCD_G0,
output LCD_G1,
output LCD_G4,
output LCD_BACKLIGHT_CTRL,
output LCD_R0,
output LCD_R1,
output UART_TX,
input UART_RX,
output I2C_SCL,
inout I2C_SDA,
input I2C_INTERRUPT,
inout SD_DAT1,
inout SD_DAT0,
output SD_CLK,
output SD_CMD,
inout SD_DAT3,
inout SD_DAT2,
output SDRAM_A0,
output SDRAM_A1,
output SDRAM_A2,
output SDRAM_A3,
output SDRAM_A4,
output SDRAM_A5,
output SDRAM_A6,
output SDRAM_A7,
output SDRAM_A8,
output SDRAM_A9,
output SDRAM_A10,
output SDRAM_A11,
output SDRAM_A12,
output SDRAM_BA0,
output SDRAM_BA1,
output SDRAM_CLK,
output SDRAM_CKE,
output SDRAM_RAS_n,
output SDRAM_CAS_n,
output SDRAM_WE_n,
output SDRAM_CE_n,
inout SDRAM_DQ0,
inout SDRAM_DQ1,
inout SDRAM_DQ2,
inout SDRAM_DQ3,
inout SDRAM_DQ4,
inout SDRAM_DQ5,
inout SDRAM_DQ6,
inout SDRAM_DQ7,
inout SDRAM_DQ8,
inout SDRAM_DQ9,
inout SDRAM_DQ10,
inout SDRAM_DQ11,
inout SDRAM_DQ12,
inout SDRAM_DQ13,
inout SDRAM_DQ14,
inout SDRAM_DQ15,
output SDRAM_DQM0,
output SDRAM_DQM1
